
module	Top_Random_Maze	(	
					input	logic clk,
					input	logic resetN,
					input	logic [10:0] pixelX, // current VGA pixel 
					input	logic [10:0] pixelY,
					input	logic startOfFrame, // short pulse every start of frame 30Hz 
					input	logic [2:0] level,
					input	logic draw_random, 
					input	logic empty_map, // empty map - when you get a surprise/win/lose

					output	logic [7:0] RGBout, // optional color output for mux 
					output	logic mazeDrawingRequest
);

parameter int MAPS_IN_LVL_NUM = 3;
parameter int LEVEL_NUM = 5;
parameter int BLOCK_ROWS = 15; //the number of rows and columns of blocks in the matrix
parameter int BLOCK_COLS = 20;

// this is the devider used to acess the right pixel 
parameter int OBJECT_NUMBER_OF_Y_BITS = 5;  // 2^5 = 32 
parameter int OBJECT_NUMBER_OF_X_BITS = 5;  // 2^5 = 32 

//the variables that are used in order to determine the current row and column
logic [BLOCK_ROWS-1:0]i; //row index
assign i = pixelY >> OBJECT_NUMBER_OF_Y_BITS;  
logic [BLOCK_COLS-1:0]j; //column index
assign j = pixelX >> OBJECT_NUMBER_OF_X_BITS;  

localparam int OBJECT_HEIGHT_Y = 1 <<  OBJECT_NUMBER_OF_Y_BITS ;
localparam int OBJECT_WIDTH_X = 1 <<  OBJECT_NUMBER_OF_X_BITS;

logic block_req_in;
logic [10:0] offsetX_in;
logic [10:0] offsetY_in;
logic [1:0] random_in;
logic [0:OBJECT_HEIGHT_Y-1][0:OBJECT_WIDTH_X-1] [8-1:0] block_object_colors_in;


bit [0:LEVEL_NUM-1] [0:MAPS_IN_LVL_NUM-1] [0:BLOCK_ROWS-1] [0:BLOCK_COLS-1] maze_bitmap  = { //[current level][random map][requested row][requested col]

{
{20'b	11111111111111111111,
20'b	11000000110000000011,
20'b	10000000011000000001,
20'b	10000000000110000001,
20'b	10000000000001100001,
20'b	10000000000000100001,
20'b	10000111111000000001,
20'b	11111100000000000001,
20'b	10000000000011000001,
20'b	10000000001100000001,
20'b	10000000111000000001,
20'b	10000000011111110001,
20'b	10000000000000010001,
20'b	10000011111100000001,
20'b	11111111111111111111},
																	
{20'b	11111111111111111111,
20'b	11000000000000000101,
20'b	11000000000001111001,
20'b	11110000000011000001,
20'b	10001100000000000001,
20'b	10000111000000000001,
20'b	10000000110000000001,
20'b	10000000000000011111,
20'b	10000000000000000001,
20'b	10000001111000000001,
20'b	11111111000000000001,
20'b	10000001110000000001,
20'b	10000000000000000001,
20'b	10000000001110000001,
20'b	11111111111111111111},

{20'b	11111111111111111111,
20'b	11000000000000000111,
20'b	10000001111100000001,
20'b	10000000001111000001,
20'b	10000000111000000001,
20'b	10000000000000000001,
20'b	10000000000000000001,
20'b	10001111100011100001,
20'b	10000000111110000001,
20'b	10000000000000000001,
20'b	10000000000000000001,
20'b	10000000000110000001,
20'b	10000000011110000001,
20'b	10000011111111110001,
20'b	11111111111111111111},
},

{
{20'b	11111111111111111111,
20'b	10100000000000000011,
20'b	10111110000000000001,
20'b	10000011110000001111,
20'b	10000000011000000001,
20'b	10000000001000000001,
20'b	10000000011000001111,
20'b	10000000110000000001,
20'b	10000011100000000001,
20'b	10000111000000000001,
20'b	10011100000000000001,
20'b	10000000000011100001,
20'b	10000000011111000001,
20'b	10000011111110000001,
20'b	11111111111111111111},
																	
{20'b	11111111111111111111,
20'b	10100000000000000101,
20'b	10100000110000000001,
20'b	10110111100000111111,
20'b	10011110000000100001,
20'b	10000011000000100001,
20'b	10000000000001100001,
20'b	10000000000011000001,
20'b	11110000000000000001,
20'b	10011000011000001111,
20'b	10001100000000001001,
20'b	10000111100000001001,
20'b	10000000111000000001,
20'b	10000000000000000001,
20'b	11111111111111111111},

{20'b	11111111111111111111,
20'b	10100000000000000111,
20'b	10011100000000000001,
20'b	10000111000000110001,
20'b	10000011000000010001,
20'b	10000011110000011001,
20'b	10000000011000001001,
20'b	10000000000000001001,
20'b	10000000000000000001,
20'b	11000111110000000001,
20'b	10100001111111000001,
20'b	10000001100000000001,
20'b	10000000111000010001,
20'b	10000111100000110001,
20'b	11111111111111111111},
},

{
{20'b	11111111111111111111,
20'b	11100000000000000011,
20'b	11111000000000001111,
20'b	10001111000001110001,
20'b	10000000000011100001,
20'b	10000000011001100001,
20'b	10001111000000110001,
20'b	10011110000000011001,
20'b	10111000000000001101,
20'b	10101100110000111101,
20'b	10100000000000000001,
20'b	10110000001111000001,
20'b	10011111000000000001,
20'b	10000000000111000001,
20'b	11111111111111111111},
																	
{20'b	11111111111111111111,
20'b	11100000000000000101,
20'b	11100011000000000001,
20'b	10100110000000000001,
20'b	10011111100000110001,
20'b	10000000000000100001,
20'b	10000000000111100001,
20'b	10000000001000000001,
20'b	10000001110000000001,
20'b	10000110000011000001,
20'b	10000000000110000001,
20'b	10000011111100010001,
20'b	10000000011111110001,
20'b	11000000000000000001,
20'b	11111111111111111111},

{20'b	11111111111111111111,
20'b	11100000000000000111,
20'b	10000000000011100001,
20'b	10000000001110000001,
20'b	10000111110000000001,
20'b	10000000111111111001,
20'b	10111111111000000001,
20'b	10000000000001100001,
20'b	10000011100000000001,
20'b	10000001111000000001,
20'b	10000110000000001001,
20'b	10000001110000001001,
20'b	10000001111100010001,
20'b	11111000000000010001,
20'b	11111111111111111111},
},

{
{20'b	11111111111111111111,
20'b	10010000001110000011,
20'b	10001111000011110001,
20'b	10000000001111000001,
20'b	10000110000000001101,
20'b	10100001110110000001,
20'b	10110000000111000001,
20'b	11110000111111111001,
20'b	10000000000011000001,
20'b	10001110110011000001,
20'b	10000110010000011101,
20'b	10000000011000000101,
20'b	10000110000111000001,
20'b	10011100001111100001,
20'b	11111111111111111111},
																	
{20'b	11111111111111111111,
20'b	10010000000000000101,
20'b	10000011111111100001,
20'b	10000000000011100001,
20'b	10000111000010000001,
20'b	10000001110110000001,
20'b	10000000000000011001,
20'b	10000000011100111001,
20'b	10011000000011000001,
20'b	10000010110011010001,
20'b	10000111110000000001,
20'b	10000000011111000001,
20'b	10000000000111000001,
20'b	10011100000001110001,
20'b	11111111111111111111},

{20'b	11111111111111111111,
20'b	10010001110000000111,
20'b	10010011000011111001,
20'b	10000000000111111001,
20'b	10011110001111000001,
20'b	10001111000000000001,
20'b	10000011100100001001,
20'b	10000000000100011001,
20'b	10000000011000010001,
20'b	10000111110001110001,
20'b	10000000111000000001,
20'b	10000000100001111001,
20'b	10001101111001111001,
20'b	10000111111000111001,
20'b	11111111111111111111},
},

{
{20'b	11111111111111111111,
20'b	11010000000000000011,
20'b	11011111110000000001,
20'b	10000100011100000001,
20'b	10000000001111010001,
20'b	10110010000010001001,
20'b	10000010000000001001,
20'b	10000110000001001001,
20'b	10001110000001000111,
20'b	10111000000111100001,
20'b	10100000011110001001,
20'b	10111001110000011001,
20'b	10011111100000111001,
20'b	10000000000011100001,
20'b	11111111111111111111},
																	
{20'b	11111111111111111111,
20'b	11010000000000000101,
20'b	10011111110000000001,
20'b	10000000111111111001,
20'b	10000000000011111101,
20'b	10000111111111000001,
20'b	10001111000001000001,
20'b	10011000000000001001,
20'b	10010000111000110001,
20'b	10011000000001110001,
20'b	10001110011111000001,
20'b	10000011110000000001,
20'b	10001110011111001001,
20'b	10000000000000001101,
20'b	11111111111111111111},

{20'b	11111111111111111111,
20'b	11010000000000000111,
20'b	10010011100000000001,
20'b	10110011110000011111,
20'b	10011000011110000001,
20'b	10000000001111100011,
20'b	10000001111110000111,
20'b	10001111110000000001,
20'b	10000000111111111001,
20'b	10011111111110000001,
20'b	10000000111000010001,
20'b	10000000011100100001,
20'b	10011110000011100001,
20'b	10000111110000000101,
20'b	11111111111111111111},
},
};

bit [0:BLOCK_ROWS-1] [0:BLOCK_COLS-1] empty_bitmap  = { //empty map - when the player wins/loses/receives a surprise

20'b	11111111111111111111,
20'b	10000000000000000001,
20'b	10000000000000000001,
20'b	10000000000000000001,
20'b	10000000000000000001,
20'b	10000000000000000001,
20'b	10000000000000000001,
20'b	10000000000000000001,
20'b	10000000000000000001,
20'b	10000000000000000001,
20'b	10000000000000000001,
20'b	10000000000000000001,
20'b	10000000000000000001,
20'b	10000000000000000001,
20'b	11111111111111111111
};

		blockBitMap blockBitMap(.block_object_colors(block_object_colors_in));

				square_object #(.OBJECT_WIDTH_X(OBJECT_WIDTH_X), .OBJECT_HEIGHT_Y(OBJECT_HEIGHT_Y)) square_object (
					.clk(clk),
					.resetN(resetN),
					.pixelX(pixelX),
					.pixelY(pixelY),
					.topLeftX(j * OBJECT_WIDTH_X), //the actual location of the TopLeft of the block
					.topLeftY(i * OBJECT_HEIGHT_Y), //the actual location of the TopLeft of the block
					.offsetX(offsetX_in),
					.offsetY(offsetY_in),
					.drawingRequest(block_req_in),
					.RGBout()
				);
				
				random #(.SIZE_BITS(2), .MIN_VAL(0), .MAX_VAL(MAPS_IN_LVL_NUM-1), .shift_num(0)) random (
					.clk(clk),
					.resetN(resetN),					
					.rise(draw_random),
					.dout(random_in)
				);	
					
				blockDraw Draw (
					.clk(clk),					
					.resetN(resetN),
					.offsetX(offsetX_in),
					.offsetY(offsetY_in),
					.InsideRectangle(block_req_in),
					.block_object_colors(block_object_colors_in),
					//if the empty_map is enabled, choose the empty bitmap. else, choose a random map from the current level
					.enable_block((empty_map) ? empty_bitmap[i][j]: maze_bitmap[level-1][random_in][i][j]), 
					.drawingRequest(mazeDrawingRequest),
					.RGBout(RGBout)
				);


endmodule 